module main;
initial $hello(1);
endmodule